
import ClientServer::*;
import FIFO::*;
import GetPut::*;

import FixedPoint::*;
import Vector::*;

import ComplexMP::*;


typedef Server#(
    Vector#(nbins, ComplexMP#(isize, fsize, psize)),
    Vector#(nbins, ComplexMP#(isize, fsize, psize))
) PitchAdjust#(numeric type nbins, numeric type isize, numeric type fsize, numeric type psize);


// s - the amount each window is shifted from the previous window.
//
// factor - the amount to adjust the pitch.
//  1.0 makes no change. 2.0 goes up an octave, 0.5 goes down an octave, etc...
module mkPitchAdjust(Integer s, FixedPoint#(isize, fsize) factor, PitchAdjust#(nbins, isize, fsize, psize) ifc) provisos(RealLiteral#(FixedPoint#(isize, fsize)));
    Vector#(nbins, Reg#(ComplexMP#(isize, fsize, psize))) inphases <- replicateM(mkRegU());
    Vector#(nbins, Reg#(ComplexMP#(isize, fsize, psize))) outphases <- replicateM(mkReg(cmplxmp(0.0, 0)));

endmodule

